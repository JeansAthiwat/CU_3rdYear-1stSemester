`timescale 1ns / 1ps

module squarewave_rom( //8x64 tile size with square pattern 
	input clk,
	input[7:0] addr, //7:6 for square-wave pattern , 5:0 for column address of that pattern
	output reg[7:0] data
    );
	 reg[7:0] addr_q;
	 always @(posedge clk) addr_q<=addr;
	 
	 always @* begin
		 case(addr_q)
		
				//0->0				
				{2'b00 , 6'd	0	}: data= 8'b	00000000	;
				{2'b00 , 6'd	1	}: data= 8'b	00000000	;
				{2'b00 , 6'd	2	}: data= 8'b	00000000	;
				{2'b00 , 6'd	3	}: data= 8'b	00000000	;
				{2'b00 , 6'd	4	}: data= 8'b	00000000	;
				{2'b00 , 6'd	5	}: data= 8'b	00000000	;
				{2'b00 , 6'd	6	}: data= 8'b	00000000	;
				{2'b00 , 6'd	7	}: data= 8'b	00000000	;
				{2'b00 , 6'd	8	}: data= 8'b	00000000	;
				{2'b00 , 6'd	9	}: data= 8'b	00000000	;
				{2'b00 , 6'd	10	}: data= 8'b	00000000	;
				{2'b00 , 6'd	11	}: data= 8'b	00000000	;
				{2'b00 , 6'd	12	}: data= 8'b	00000000	;
				{2'b00 , 6'd	13	}: data= 8'b	00000000	;
				{2'b00 , 6'd	14	}: data= 8'b	00000000	;
				{2'b00 , 6'd	15	}: data= 8'b	00000000	;
				{2'b00 , 6'd	16	}: data= 8'b	00000000	;
				{2'b00 , 6'd	17	}: data= 8'b	00000000	;
				{2'b00 , 6'd	18	}: data= 8'b	00000000	;
				{2'b00 , 6'd	19	}: data= 8'b	00000000	;
				{2'b00 , 6'd	20	}: data= 8'b	00000000	;
				{2'b00 , 6'd	21	}: data= 8'b	00000000	;
				{2'b00 , 6'd	22	}: data= 8'b	00000000	;
				{2'b00 , 6'd	23	}: data= 8'b	00000000	;
				{2'b00 , 6'd	24	}: data= 8'b	00000000	;
				{2'b00 , 6'd	25	}: data= 8'b	00000000	;
				{2'b00 , 6'd	26	}: data= 8'b	00000000	;
				{2'b00 , 6'd	27	}: data= 8'b	00000000	;
				{2'b00 , 6'd	28	}: data= 8'b	00000000	;
				{2'b00 , 6'd	29	}: data= 8'b	00000000	;
				{2'b00 , 6'd	30	}: data= 8'b	00000000	;
				{2'b00 , 6'd	31	}: data= 8'b	00000000	;
				{2'b00 , 6'd	32	}: data= 8'b	00000000	;
				{2'b00 , 6'd	33	}: data= 8'b	00000000	;
				{2'b00 , 6'd	34	}: data= 8'b	00000000	;
				{2'b00 , 6'd	35	}: data= 8'b	00000000	;
				{2'b00 , 6'd	36	}: data= 8'b	00000000	;
				{2'b00 , 6'd	37	}: data= 8'b	00000000	;
				{2'b00 , 6'd	38	}: data= 8'b	00000000	;
				{2'b00 , 6'd	39	}: data= 8'b	00000000	;
				{2'b00 , 6'd	40	}: data= 8'b	00000000	;
				{2'b00 , 6'd	41	}: data= 8'b	00000000	;
				{2'b00 , 6'd	42	}: data= 8'b	00000000	;
				{2'b00 , 6'd	43	}: data= 8'b	00000000	;
				{2'b00 , 6'd	44	}: data= 8'b	00000000	;
				{2'b00 , 6'd	45	}: data= 8'b	00000000	;
				{2'b00 , 6'd	46	}: data= 8'b	00000000	;
				{2'b00 , 6'd	47	}: data= 8'b	00000000	;
				{2'b00 , 6'd	48	}: data= 8'b	00000000	;
				{2'b00 , 6'd	49	}: data= 8'b	00000000	;
				{2'b00 , 6'd	50	}: data= 8'b	00000000	;
				{2'b00 , 6'd	51	}: data= 8'b	00000000	;
				{2'b00 , 6'd	52	}: data= 8'b	00000000	;
				{2'b00 , 6'd	53	}: data= 8'b	00000000	;
				{2'b00 , 6'd	54	}: data= 8'b	00000000	;
				{2'b00 , 6'd	55	}: data= 8'b	00000000	;
				{2'b00 , 6'd	56	}: data= 8'b	00000000	;
				{2'b00 , 6'd	57	}: data= 8'b	00000000	;
				{2'b00 , 6'd	58	}: data= 8'b	00000000	;
				{2'b00 , 6'd	59	}: data= 8'b	00000000	;
				{2'b00 , 6'd	60	}: data= 8'b	00000000	;
				{2'b00 , 6'd	61	}: data= 8'b	00000000	;
				{2'b00 , 6'd	62	}: data= 8'b	00000000	;
				{2'b00 , 6'd	63	}: data= 8'b	11111111	;
								
				//0->1				
				{2'b01, 6'd	0	}: data= 8'b	00001111	;
				{2'b01, 6'd	1	}: data= 8'b	00001000	;
				{2'b01, 6'd	2	}: data= 8'b	00001000	;
				{2'b01, 6'd	3	}: data= 8'b	00001000	;
				{2'b01, 6'd	4	}: data= 8'b	00001000	;
				{2'b01, 6'd	5	}: data= 8'b	00001000	;
				{2'b01, 6'd	6	}: data= 8'b	00001000	;
				{2'b01, 6'd	7	}: data= 8'b	00001000	;
				{2'b01, 6'd	8	}: data= 8'b	00001000	;
				{2'b01, 6'd	9	}: data= 8'b	00001000	;
				{2'b01, 6'd	10	}: data= 8'b	00001000	;
				{2'b01, 6'd	11	}: data= 8'b	00001000	;
				{2'b01, 6'd	12	}: data= 8'b	00001000	;
				{2'b01, 6'd	13	}: data= 8'b	00001000	;
				{2'b01, 6'd	14	}: data= 8'b	00001000	;
				{2'b01, 6'd	15	}: data= 8'b	00001000	;
				{2'b01, 6'd	16	}: data= 8'b	00001000	;
				{2'b01, 6'd	17	}: data= 8'b	00001000	;
				{2'b01, 6'd	18	}: data= 8'b	00001000	;
				{2'b01, 6'd	19	}: data= 8'b	00001000	;
				{2'b01, 6'd	20	}: data= 8'b	00001000	;
				{2'b01, 6'd	21	}: data= 8'b	00001000	;
				{2'b01, 6'd	22	}: data= 8'b	00001000	;
				{2'b01, 6'd	23	}: data= 8'b	00001000	;
				{2'b01, 6'd	24	}: data= 8'b	00001000	;
				{2'b01, 6'd	25	}: data= 8'b	00001000	;
				{2'b01, 6'd	26	}: data= 8'b	00001000	;
				{2'b01, 6'd	27	}: data= 8'b	00001000	;
				{2'b01, 6'd	28	}: data= 8'b	00001000	;
				{2'b01, 6'd	29	}: data= 8'b	00001000	;
				{2'b01, 6'd	30	}: data= 8'b	00001000	;
				{2'b01, 6'd	31	}: data= 8'b	00001000	;
				{2'b01, 6'd	32	}: data= 8'b	00001000	;
				{2'b01, 6'd	33	}: data= 8'b	00001000	;
				{2'b01, 6'd	34	}: data= 8'b	00001000	;
				{2'b01, 6'd	35	}: data= 8'b	00001000	;
				{2'b01, 6'd	36	}: data= 8'b	00001000	;
				{2'b01, 6'd	37	}: data= 8'b	00001000	;
				{2'b01, 6'd	38	}: data= 8'b	00001000	;
				{2'b01, 6'd	39	}: data= 8'b	00001000	;
				{2'b01, 6'd	40	}: data= 8'b	00001000	;
				{2'b01, 6'd	41	}: data= 8'b	00001000	;
				{2'b01, 6'd	42	}: data= 8'b	00001000	;
				{2'b01, 6'd	43	}: data= 8'b	00001000	;
				{2'b01, 6'd	44	}: data= 8'b	00001000	;
				{2'b01, 6'd	45	}: data= 8'b	00001000	;
				{2'b01, 6'd	46	}: data= 8'b	00001000	;
				{2'b01, 6'd	47	}: data= 8'b	00001000	;
				{2'b01, 6'd	48	}: data= 8'b	00001000	;
				{2'b01, 6'd	49	}: data= 8'b	00001000	;
				{2'b01, 6'd	50	}: data= 8'b	00001000	;
				{2'b01, 6'd	51	}: data= 8'b	00001000	;
				{2'b01, 6'd	52	}: data= 8'b	00001000	;
				{2'b01, 6'd	53	}: data= 8'b	00001000	;
				{2'b01, 6'd	54	}: data= 8'b	00001000	;
				{2'b01, 6'd	55	}: data= 8'b	00001000	;
				{2'b01, 6'd	56	}: data= 8'b	00001000	;
				{2'b01, 6'd	57	}: data= 8'b	00001000	;
				{2'b01, 6'd	58	}: data= 8'b	00001000	;
				{2'b01, 6'd	59	}: data= 8'b	00001000	;
				{2'b01, 6'd	60	}: data= 8'b	00001000	;
				{2'b01, 6'd	61	}: data= 8'b	00001000	;
				{2'b01, 6'd	62	}: data= 8'b	00001000	;
				{2'b01, 6'd	63	}: data= 8'b	11111000	;
								
								
				//1->1				
				{2'b11 , 6'd	0	}: data= 8'b	11111111	;
				{2'b11 , 6'd	1	}: data= 8'b	00000000	;
				{2'b11 , 6'd	2	}: data= 8'b	00000000	;
				{2'b11 , 6'd	3	}: data= 8'b	00000000	;
				{2'b11 , 6'd	4	}: data= 8'b	00000000	;
				{2'b11 , 6'd	5	}: data= 8'b	00000000	;
				{2'b11 , 6'd	6	}: data= 8'b	00000000	;
				{2'b11 , 6'd	7	}: data= 8'b	00000000	;
				{2'b11 , 6'd	8	}: data= 8'b	00000000	;
				{2'b11 , 6'd	9	}: data= 8'b	00000000	;
				{2'b11 , 6'd	10	}: data= 8'b	00000000	;
				{2'b11 , 6'd	11	}: data= 8'b	00000000	;
				{2'b11 , 6'd	12	}: data= 8'b	00000000	;
				{2'b11 , 6'd	13	}: data= 8'b	00000000	;
				{2'b11 , 6'd	14	}: data= 8'b	00000000	;
				{2'b11 , 6'd	15	}: data= 8'b	00000000	;
				{2'b11 , 6'd	16	}: data= 8'b	00000000	;
				{2'b11 , 6'd	17	}: data= 8'b	00000000	;
				{2'b11 , 6'd	18	}: data= 8'b	00000000	;
				{2'b11 , 6'd	19	}: data= 8'b	00000000	;
				{2'b11 , 6'd	20	}: data= 8'b	00000000	;
				{2'b11 , 6'd	21	}: data= 8'b	00000000	;
				{2'b11 , 6'd	22	}: data= 8'b	00000000	;
				{2'b11 , 6'd	23	}: data= 8'b	00000000	;
				{2'b11 , 6'd	24	}: data= 8'b	00000000	;
				{2'b11 , 6'd	25	}: data= 8'b	00000000	;
				{2'b11 , 6'd	26	}: data= 8'b	00000000	;
				{2'b11 , 6'd	27	}: data= 8'b	00000000	;
				{2'b11 , 6'd	28	}: data= 8'b	00000000	;
				{2'b11 , 6'd	29	}: data= 8'b	00000000	;
				{2'b11 , 6'd	30	}: data= 8'b	00000000	;
				{2'b11 , 6'd	31	}: data= 8'b	00000000	;
				{2'b11 , 6'd	32	}: data= 8'b	00000000	;
				{2'b11 , 6'd	33	}: data= 8'b	00000000	;
				{2'b11 , 6'd	34	}: data= 8'b	00000000	;
				{2'b11 , 6'd	35	}: data= 8'b	00000000	;
				{2'b11 , 6'd	36	}: data= 8'b	00000000	;
				{2'b11 , 6'd	37	}: data= 8'b	00000000	;
				{2'b11 , 6'd	38	}: data= 8'b	00000000	;
				{2'b11 , 6'd	39	}: data= 8'b	00000000	;
				{2'b11 , 6'd	40	}: data= 8'b	00000000	;
				{2'b11 , 6'd	41	}: data= 8'b	00000000	;
				{2'b11 , 6'd	42	}: data= 8'b	00000000	;
				{2'b11 , 6'd	43	}: data= 8'b	00000000	;
				{2'b11 , 6'd	44	}: data= 8'b	00000000	;
				{2'b11 , 6'd	45	}: data= 8'b	00000000	;
				{2'b11 , 6'd	46	}: data= 8'b	00000000	;
				{2'b11 , 6'd	47	}: data= 8'b	00000000	;
				{2'b11 , 6'd	48	}: data= 8'b	00000000	;
				{2'b11 , 6'd	49	}: data= 8'b	00000000	;
				{2'b11 , 6'd	50	}: data= 8'b	00000000	;
				{2'b11 , 6'd	51	}: data= 8'b	00000000	;
				{2'b11 , 6'd	52	}: data= 8'b	00000000	;
				{2'b11 , 6'd	53	}: data= 8'b	00000000	;
				{2'b11 , 6'd	54	}: data= 8'b	00000000	;
				{2'b11 , 6'd	55	}: data= 8'b	00000000	;
				{2'b11 , 6'd	56	}: data= 8'b	00000000	;
				{2'b11 , 6'd	57	}: data= 8'b	00000000	;
				{2'b11 , 6'd	58	}: data= 8'b	00000000	;
				{2'b11 , 6'd	59	}: data= 8'b	00000000	;
				{2'b11 , 6'd	60	}: data= 8'b	00000000	;
				{2'b11 , 6'd	61	}: data= 8'b	00000000	;
				{2'b11 , 6'd	62	}: data= 8'b	00000000	;
				{2'b11 , 6'd	63	}: data= 8'b	00000000	;
								
								
				//1->0				
				{2'b10 , 6'd	0	}: data= 8'b	11110000	;
				{2'b10 , 6'd	1	}: data= 8'b	00010000	;
				{2'b10 , 6'd	2	}: data= 8'b	00010000	;
				{2'b10 , 6'd	3	}: data= 8'b	00010000	;
				{2'b10 , 6'd	4	}: data= 8'b	00010000	;
				{2'b10 , 6'd	5	}: data= 8'b	00010000	;
				{2'b10 , 6'd	6	}: data= 8'b	00010000	;
				{2'b10 , 6'd	7	}: data= 8'b	00010000	;
				{2'b10 , 6'd	8	}: data= 8'b	00010000	;
				{2'b10 , 6'd	9	}: data= 8'b	00010000	;
				{2'b10 , 6'd	10	}: data= 8'b	00010000	;
				{2'b10 , 6'd	11	}: data= 8'b	00010000	;
				{2'b10 , 6'd	12	}: data= 8'b	00010000	;
				{2'b10 , 6'd	13	}: data= 8'b	00010000	;
				{2'b10 , 6'd	14	}: data= 8'b	00010000	;
				{2'b10 , 6'd	15	}: data= 8'b	00010000	;
				{2'b10 , 6'd	16	}: data= 8'b	00010000	;
				{2'b10 , 6'd	17	}: data= 8'b	00010000	;
				{2'b10 , 6'd	18	}: data= 8'b	00010000	;
				{2'b10 , 6'd	19	}: data= 8'b	00010000	;
				{2'b10 , 6'd	20	}: data= 8'b	00010000	;
				{2'b10 , 6'd	21	}: data= 8'b	00010000	;
				{2'b10 , 6'd	22	}: data= 8'b	00010000	;
				{2'b10 , 6'd	23	}: data= 8'b	00010000	;
				{2'b10 , 6'd	24	}: data= 8'b	00010000	;
				{2'b10 , 6'd	25	}: data= 8'b	00010000	;
				{2'b10 , 6'd	26	}: data= 8'b	00010000	;
				{2'b10 , 6'd	27	}: data= 8'b	00010000	;
				{2'b10 , 6'd	28	}: data= 8'b	00010000	;
				{2'b10 , 6'd	29	}: data= 8'b	00010000	;
				{2'b10 , 6'd	30	}: data= 8'b	00010000	;
				{2'b10 , 6'd	31	}: data= 8'b	00010000	;
				{2'b10 , 6'd	32	}: data= 8'b	00010000	;
				{2'b10 , 6'd	33	}: data= 8'b	00010000	;
				{2'b10 , 6'd	34	}: data= 8'b	00010000	;
				{2'b10 , 6'd	35	}: data= 8'b	00010000	;
				{2'b10 , 6'd	36	}: data= 8'b	00010000	;
				{2'b10 , 6'd	37	}: data= 8'b	00010000	;
				{2'b10 , 6'd	38	}: data= 8'b	00010000	;
				{2'b10 , 6'd	39	}: data= 8'b	00010000	;
				{2'b10 , 6'd	40	}: data= 8'b	00010000	;
				{2'b10 , 6'd	41	}: data= 8'b	00010000	;
				{2'b10 , 6'd	42	}: data= 8'b	00010000	;
				{2'b10 , 6'd	43	}: data= 8'b	00010000	;
				{2'b10 , 6'd	44	}: data= 8'b	00010000	;
				{2'b10 , 6'd	45	}: data= 8'b	00010000	;
				{2'b10 , 6'd	46	}: data= 8'b	00010000	;
				{2'b10 , 6'd	47	}: data= 8'b	00010000	;
				{2'b10 , 6'd	48	}: data= 8'b	00010000	;
				{2'b10 , 6'd	49	}: data= 8'b	00010000	;
				{2'b10 , 6'd	50	}: data= 8'b	00010000	;
				{2'b10 , 6'd	51	}: data= 8'b	00010000	;
				{2'b10 , 6'd	52	}: data= 8'b	00010000	;
				{2'b10 , 6'd	53	}: data= 8'b	00010000	;
				{2'b10 , 6'd	54	}: data= 8'b	00010000	;
				{2'b10 , 6'd	55	}: data= 8'b	00010000	;
				{2'b10 , 6'd	56	}: data= 8'b	00010000	;
				{2'b10 , 6'd	57	}: data= 8'b	00010000	;
				{2'b10 , 6'd	58	}: data= 8'b	00010000	;
				{2'b10 , 6'd	59	}: data= 8'b	00010000	;
				{2'b10 , 6'd	60	}: data= 8'b	00010000	;
				{2'b10 , 6'd	61	}: data= 8'b	00010000	;
				{2'b10 , 6'd	62	}: data= 8'b	00010000	;
				{2'b10 , 6'd	63	}: data= 8'b	00011111	;

		 
		 
		 endcase
	end


endmodule
